module LA_MUX #(parameter pADDR_WIDTH = 12,
                parameter pDATA_WIDTH = 32)
(
	input wire ALCLK,
	input wire ARESET_N,
	input wire [0:0] USER_PRJ_SEL,
	input wire [63:0] la_data,
	input wire [63:0] la_data,
	input wire [63:0] la_data,
	input wire [63:0] la_data
	output wire [63:0] la_data
);

endmodule //LA_MUX

