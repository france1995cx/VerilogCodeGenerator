module USER_SUB_SYS #(parameter pADDR_WIDTH = 12,
                      parameter pDATA_WIDTH = 32)
(
	input wire [pADDR_WIDTH-1:0] a_ls_araddr,
	input wire a_ls_arvalid,
	input wire [pADDR_WIDTH-1:0] a_ls_awaddr,
	input wire a_ls_awvalid,
	input wire [pDATA_WIDTH-1:0] a_ls_wdata,
	input wire a_ls_wstrb,
	input wire a_ls_wvalid,
	input wire a_lsrready,
	input wire a_sm_tready,
	input wire [pDATA_WIDTH-1:0] a_ss_tdata,
	input wire [2:0] a_ss_tid,
	input wire a_ss_tkeep,
	input wire a_ss_tlast,
	input wire [3:0] a_ss_tstrb,
	input wire a_ss_tvalid
	output wire a_ls_arready,
	output wire a_ls_awready,
	output wire [pDATA_WIDTH-1:0] a_ls_rdata,
	output wire a_ls_rvalid,
	output wire a_ls_wready,
	output wire [pDATA_WIDTH-1:0] a_sm_tdata,
	output wire [2:0] a_sm_tid,
	output wire a_sm_tkeep,
	output wire a_sm_tlast,
	output wire [3:0] a_sm_tstrb,
	output wire a_sm_tvalid,
	output wire a_ss_tready,
	output wire hi_pri_req,
	output wire [63:0] la_data,
	output wire user_irq
);
wire ALCLK;
wire ARESET_N;
wire [0:0] USER_PRJ_SEL;
wire [pADDR_WIDTH-1:0] a_ls_araddr;
wire a_ls_arvalid;
wire [pADDR_WIDTH-1:0] a_ls_awaddr;
wire a_ls_awvalid;
wire [pDATA_WIDTH-1:0] a_ls_wdata;
wire a_ls_wstrb;
wire a_ls_wvalid;
wire a_lsrready;
wire arready;
wire arready;
wire arready;
wire arready;
wire awready;
wire awready;
wire awready;
wire awready;
wire [pDATA_WIDTH-1:0] rdata;
wire [pDATA_WIDTH-1:0] rdata;
wire [pDATA_WIDTH-1:0] rdata;
wire [pDATA_WIDTH-1:0] rdata;
wire rvalid;
wire rvalid;
wire rvalid;
wire rvalid;
wire wready;
wire wready;
wire wready;
wire wreadywire Arvalid_0;
wire [pDATA_WIDTH-1:0] Wdata;
wire [pDATA_WIDTH-1:0] Wdata;
wire [pDATA_WIDTH-1:0] Wdata;
wire [pDATA_WIDTH-1:0] Wdata;
wire a_ls_arready;
wire a_ls_awready;
wire [pDATA_WIDTH-1:0] a_ls_rdata;
wire a_ls_rvalid;
wire a_ls_wready;
wire [pADDR_WIDTH-1:0] araddr;
wire [pADDR_WIDTH-1:0] araddr;
wire [pADDR_WIDTH-1:0] araddr;
wire [pADDR_WIDTH-1:0] araddr;
wire arvalid_1;
wire arvalid_2;
wire arvalid_3;
wire [pADDR_WIDTH-1:0] awaddr;
wire [pADDR_WIDTH-1:0] awaddr;
wire [pADDR_WIDTH-1:0] awaddr;
wire [pADDR_WIDTH-1:0] awaddr;
wire awvalid_0;
wire awvalid_1;
wire awvalid_2;
wire awvalid_3;
wire rready;
wire rready;
wire rready;
wire rready;
wire wstrb_0;
wire wstrb_1;
wire wstrb_2;
wire wstrb_3;
wire wvalid_0;
wire wvalid_1;
wire wvalid_2;
wire wvalid_3
AXIL_SLAV #(.pADDR_WIDTH(12),
            .pDATA_WIDTH(32))AXIL_SLAV (
                                     .ALCLK (ALCLK).
                                     .ARESET_N (ARESET_N).
                                     .USER_PRJ_SEL (USER_PRJ_SEL).
                                     .a_ls_araddr (a_ls_araddr).
                                     .a_ls_arvalid (a_ls_arvalid).
                                     .a_ls_awaddr (a_ls_awaddr).
                                     .a_ls_awvalid (a_ls_awvalid).
                                     .a_ls_wdata (a_ls_wdata).
                                     .a_ls_wstrb (a_ls_wstrb).
                                     .a_ls_wvalid (a_ls_wvalid).
                                     .a_lsrready (a_lsrready).
                                     .arready (arready).
                                     .arready (arready).
                                     .arready (arready).
                                     .arready (arready).
                                     .awready (awready).
                                     .awready (awready).
                                     .awready (awready).
                                     .awready (awready).
                                     .rdata (rdata).
                                     .rdata (rdata).
                                     .rdata (rdata).
                                     .rdata (rdata).
                                     .rvalid (rvalid).
                                     .rvalid (rvalid).
                                     .rvalid (rvalid).
                                     .rvalid (rvalid).
                                     .wready (wready).
                                     .wready (wready).
                                     .wready (wready).
                                     .wready (wready).
                                     .Arvalid_0 (Arvalid_0).
                                     .Wdata (Wdata).
                                     .Wdata (Wdata).
                                     .Wdata (Wdata).
                                     .Wdata (Wdata).
                                     .a_ls_arready (a_ls_arready).
                                     .a_ls_awready (a_ls_awready).
                                     .a_ls_rdata (a_ls_rdata).
                                     .a_ls_rvalid (a_ls_rvalid).
                                     .a_ls_wready (a_ls_wready).
                                     .araddr (araddr).
                                     .araddr (araddr).
                                     .araddr (araddr).
                                     .araddr (araddr).
                                     .arvalid_1 (arvalid_1).
                                     .arvalid_2 (arvalid_2).
                                     .arvalid_3 (arvalid_3).
                                     .awaddr (awaddr).
                                     .awaddr (awaddr).
                                     .awaddr (awaddr).
                                     .awaddr (awaddr).
                                     .awvalid_0 (awvalid_0).
                                     .awvalid_1 (awvalid_1).
                                     .awvalid_2 (awvalid_2).
                                     .awvalid_3 (awvalid_3).
                                     .rready (rready).
                                     .rready (rready).
                                     .rready (rready).
                                     .rready (rready).
                                     .wstrb_0 (wstrb_0).
                                     .wstrb_1 (wstrb_1).
                                     .wstrb_2 (wstrb_2).
                                     .wstrb_3 (wstrb_3).
                                     .wvalid_0 (wvalid_0).
                                     .wvalid_1 (wvalid_1).
                                     .wvalid_2 (wvalid_2).
                                     .wvalid_3 (wvalid_3).
                                     );wire ALCLK;
wire ALCLK;
wire ALCLK;
wire ALCLK;
wire ARESET_N;
wire ARESET_N;
wire ARESET_N;
wire ARESET_N;
wire ASCLK;
wire ASCLK;
wire ASCLK;
wire ASCLK;
wire Arvalid_0;
wire USER_CLK2;
wire USER_CLK2;
wire USER_CLK2;
wire USER_CLK2;
wire [pDATA_WIDTH-1:0] Wdata;
wire [pDATA_WIDTH-1:0] Wdata;
wire [pDATA_WIDTH-1:0] Wdata;
wire [pDATA_WIDTH-1:0] Wdata;
wire [pADDR_WIDTH-1:0] araddr;
wire [pADDR_WIDTH-1:0] araddr;
wire [pADDR_WIDTH-1:0] araddr;
wire [pADDR_WIDTH-1:0] araddr;
wire arvalid_1;
wire arvalid_2;
wire arvalid_3;
wire [pADDR_WIDTH-1:0] awaddr;
wire [pADDR_WIDTH-1:0] awaddr;
wire [pADDR_WIDTH-1:0] awaddr;
wire [pADDR_WIDTH-1:0] awaddr;
wire awvalid_0;
wire awvalid_1;
wire awvalid_2;
wire awvalid_3;
wire rready;
wire rready;
wire rready;
wire rready;
wire sm_tready;
wire sm_tready;
wire sm_tready;
wire sm_tready;
wire [pDATA_WIDTH-1:0] ss_tdata;
wire [pDATA_WIDTH-1:0] ss_tdata;
wire [pDATA_WIDTH-1:0] ss_tdata;
wire [pDATA_WIDTH-1:0] ss_tdata;
wire [2:0] ss_tid;
wire [2:0] ss_tid;
wire [2:0] ss_tid;
wire [2:0] ss_tid;
wire ss_tkeep;
wire ss_tkeep;
wire ss_tkeep;
wire ss_tkeep;
wire ss_tlast;
wire ss_tlast;
wire ss_tlast;
wire ss_tlast;
wire [3:0] ss_tstrb;
wire [3:0] ss_tstrb;
wire [3:0] ss_tstrb;
wire [3:0] ss_tstrb;
wire ss_tvalid_0;
wire ss_tvalid_1;
wire ss_tvalid_2;
wire ss_tvalid_3;
wire wstrb_0;
wire wstrb_1;
wire wstrb_2;
wire wstrb_3;
wire wvalid_0;
wire wvalid_1;
wire wvalid_2;
wire wvalid_3wire arready;
wire arready;
wire arready;
wire arready;
wire awready;
wire awready;
wire awready;
wire awready;
wire hi_pri_req;
wire hi_pri_req;
wire hi_pri_req;
wire hi_pri_req;
wire [63:0] la_data;
wire [63:0] la_data;
wire [63:0] la_data;
wire [63:0] la_data;
wire [pDATA_WIDTH-1:0] rdata;
wire [pDATA_WIDTH-1:0] rdata;
wire [pDATA_WIDTH-1:0] rdata;
wire [pDATA_WIDTH-1:0] rdata;
wire rvalid;
wire rvalid;
wire rvalid;
wire rvalid;
wire [pDATA_WIDTH-1:0] sm_tdata;
wire [pDATA_WIDTH-1:0] sm_tdata;
wire [pDATA_WIDTH-1:0] sm_tdata;
wire [pDATA_WIDTH-1:0] sm_tdata;
wire [2:0] sm_tid;
wire [2:0] sm_tid;
wire [2:0] sm_tid;
wire [2:0] sm_tid;
wire sm_tkeep;
wire sm_tkeep;
wire sm_tkeep;
wire sm_tkeep;
wire sm_tlast;
wire sm_tlast;
wire sm_tlast;
wire sm_tlast;
wire [3:0] sm_tstrb;
wire [3:0] sm_tstrb;
wire [3:0] sm_tstrb;
wire [3:0] sm_tstrb;
wire sm_tvalid;
wire sm_tvalid;
wire sm_tvalid;
wire sm_tvalid;
wire ss_tready;
wire ss_tready;
wire ss_tready;
wire ss_tready;
wire user_irq;
wire user_irq;
wire user_irq;
wire user_irq;
wire wready;
wire wready;
wire wready;
wire wready
USER_PRJ #(.pADDR_WIDTH(12),
           .pDATA_WIDTH(32))USER_PRJ (
                                   .ALCLK (ALCLK).
                                   .ALCLK (ALCLK).
                                   .ALCLK (ALCLK).
                                   .ALCLK (ALCLK).
                                   .ARESET_N (ARESET_N).
                                   .ARESET_N (ARESET_N).
                                   .ARESET_N (ARESET_N).
                                   .ARESET_N (ARESET_N).
                                   .ASCLK (ASCLK).
                                   .ASCLK (ASCLK).
                                   .ASCLK (ASCLK).
                                   .ASCLK (ASCLK).
                                   .Arvalid_0 (Arvalid_0).
                                   .USER_CLK2 (USER_CLK2).
                                   .USER_CLK2 (USER_CLK2).
                                   .USER_CLK2 (USER_CLK2).
                                   .USER_CLK2 (USER_CLK2).
                                   .Wdata (Wdata).
                                   .Wdata (Wdata).
                                   .Wdata (Wdata).
                                   .Wdata (Wdata).
                                   .araddr (araddr).
                                   .araddr (araddr).
                                   .araddr (araddr).
                                   .araddr (araddr).
                                   .arvalid_1 (arvalid_1).
                                   .arvalid_2 (arvalid_2).
                                   .arvalid_3 (arvalid_3).
                                   .awaddr (awaddr).
                                   .awaddr (awaddr).
                                   .awaddr (awaddr).
                                   .awaddr (awaddr).
                                   .awvalid_0 (awvalid_0).
                                   .awvalid_1 (awvalid_1).
                                   .awvalid_2 (awvalid_2).
                                   .awvalid_3 (awvalid_3).
                                   .rready (rready).
                                   .rready (rready).
                                   .rready (rready).
                                   .rready (rready).
                                   .sm_tready (sm_tready).
                                   .sm_tready (sm_tready).
                                   .sm_tready (sm_tready).
                                   .sm_tready (sm_tready).
                                   .ss_tdata (ss_tdata).
                                   .ss_tdata (ss_tdata).
                                   .ss_tdata (ss_tdata).
                                   .ss_tdata (ss_tdata).
                                   .ss_tid (ss_tid).
                                   .ss_tid (ss_tid).
                                   .ss_tid (ss_tid).
                                   .ss_tid (ss_tid).
                                   .ss_tkeep (ss_tkeep).
                                   .ss_tkeep (ss_tkeep).
                                   .ss_tkeep (ss_tkeep).
                                   .ss_tkeep (ss_tkeep).
                                   .ss_tlast (ss_tlast).
                                   .ss_tlast (ss_tlast).
                                   .ss_tlast (ss_tlast).
                                   .ss_tlast (ss_tlast).
                                   .ss_tstrb (ss_tstrb).
                                   .ss_tstrb (ss_tstrb).
                                   .ss_tstrb (ss_tstrb).
                                   .ss_tstrb (ss_tstrb).
                                   .ss_tvalid_0 (ss_tvalid_0).
                                   .ss_tvalid_1 (ss_tvalid_1).
                                   .ss_tvalid_2 (ss_tvalid_2).
                                   .ss_tvalid_3 (ss_tvalid_3).
                                   .wstrb_0 (wstrb_0).
                                   .wstrb_1 (wstrb_1).
                                   .wstrb_2 (wstrb_2).
                                   .wstrb_3 (wstrb_3).
                                   .wvalid_0 (wvalid_0).
                                   .wvalid_1 (wvalid_1).
                                   .wvalid_2 (wvalid_2).
                                   .wvalid_3 (wvalid_3).
                                   .arready (arready).
                                   .arready (arready).
                                   .arready (arready).
                                   .arready (arready).
                                   .awready (awready).
                                   .awready (awready).
                                   .awready (awready).
                                   .awready (awready).
                                   .hi_pri_req (hi_pri_req).
                                   .hi_pri_req (hi_pri_req).
                                   .hi_pri_req (hi_pri_req).
                                   .hi_pri_req (hi_pri_req).
                                   .la_data (la_data).
                                   .la_data (la_data).
                                   .la_data (la_data).
                                   .la_data (la_data).
                                   .rdata (rdata).
                                   .rdata (rdata).
                                   .rdata (rdata).
                                   .rdata (rdata).
                                   .rvalid (rvalid).
                                   .rvalid (rvalid).
                                   .rvalid (rvalid).
                                   .rvalid (rvalid).
                                   .sm_tdata (sm_tdata).
                                   .sm_tdata (sm_tdata).
                                   .sm_tdata (sm_tdata).
                                   .sm_tdata (sm_tdata).
                                   .sm_tid (sm_tid).
                                   .sm_tid (sm_tid).
                                   .sm_tid (sm_tid).
                                   .sm_tid (sm_tid).
                                   .sm_tkeep (sm_tkeep).
                                   .sm_tkeep (sm_tkeep).
                                   .sm_tkeep (sm_tkeep).
                                   .sm_tkeep (sm_tkeep).
                                   .sm_tlast (sm_tlast).
                                   .sm_tlast (sm_tlast).
                                   .sm_tlast (sm_tlast).
                                   .sm_tlast (sm_tlast).
                                   .sm_tstrb (sm_tstrb).
                                   .sm_tstrb (sm_tstrb).
                                   .sm_tstrb (sm_tstrb).
                                   .sm_tstrb (sm_tstrb).
                                   .sm_tvalid (sm_tvalid).
                                   .sm_tvalid (sm_tvalid).
                                   .sm_tvalid (sm_tvalid).
                                   .sm_tvalid (sm_tvalid).
                                   .ss_tready (ss_tready).
                                   .ss_tready (ss_tready).
                                   .ss_tready (ss_tready).
                                   .ss_tready (ss_tready).
                                   .user_irq (user_irq).
                                   .user_irq (user_irq).
                                   .user_irq (user_irq).
                                   .user_irq (user_irq).
                                   .wready (wready).
                                   .wready (wready).
                                   .wready (wready).
                                   .wready (wready).
                                   );wire ARESET_N;
wire ASCLK;
wire [0:0] USER_PRJ_SEL;
wire [pDATA_WIDTH-1:0] a_ss_tdata;
wire [2:0] a_ss_tid;
wire a_ss_tkeep;
wire a_ss_tlast;
wire [3:0] a_ss_tstrb;
wire a_ss_tvalid;
wire ss_tready;
wire ss_tready;
wire ss_tready;
wire ss_treadywire a_ss_tready;
wire [pDATA_WIDTH-1:0] ss_tdata;
wire [pDATA_WIDTH-1:0] ss_tdata;
wire [pDATA_WIDTH-1:0] ss_tdata;
wire [pDATA_WIDTH-1:0] ss_tdata;
wire [2:0] ss_tid;
wire [2:0] ss_tid;
wire [2:0] ss_tid;
wire [2:0] ss_tid;
wire ss_tkeep;
wire ss_tkeep;
wire ss_tkeep;
wire ss_tkeep;
wire ss_tlast;
wire ss_tlast;
wire ss_tlast;
wire ss_tlast;
wire [3:0] ss_tstrb;
wire [3:0] ss_tstrb;
wire [3:0] ss_tstrb;
wire [3:0] ss_tstrb;
wire ss_tvalid_0;
wire ss_tvalid_1;
wire ss_tvalid_2;
wire ss_tvalid_3
AXIS_SLAV #(.pADDR_WIDTH(12),
            .pDATA_WIDTH(32))AXIS_SLAV (
                                     .ARESET_N (ARESET_N).
                                     .ASCLK (ASCLK).
                                     .USER_PRJ_SEL (USER_PRJ_SEL).
                                     .a_ss_tdata (a_ss_tdata).
                                     .a_ss_tid (a_ss_tid).
                                     .a_ss_tkeep (a_ss_tkeep).
                                     .a_ss_tlast (a_ss_tlast).
                                     .a_ss_tstrb (a_ss_tstrb).
                                     .a_ss_tvalid (a_ss_tvalid).
                                     .ss_tready (ss_tready).
                                     .ss_tready (ss_tready).
                                     .ss_tready (ss_tready).
                                     .ss_tready (ss_tready).
                                     .a_ss_tready (a_ss_tready).
                                     .ss_tdata (ss_tdata).
                                     .ss_tdata (ss_tdata).
                                     .ss_tdata (ss_tdata).
                                     .ss_tdata (ss_tdata).
                                     .ss_tid (ss_tid).
                                     .ss_tid (ss_tid).
                                     .ss_tid (ss_tid).
                                     .ss_tid (ss_tid).
                                     .ss_tkeep (ss_tkeep).
                                     .ss_tkeep (ss_tkeep).
                                     .ss_tkeep (ss_tkeep).
                                     .ss_tkeep (ss_tkeep).
                                     .ss_tlast (ss_tlast).
                                     .ss_tlast (ss_tlast).
                                     .ss_tlast (ss_tlast).
                                     .ss_tlast (ss_tlast).
                                     .ss_tstrb (ss_tstrb).
                                     .ss_tstrb (ss_tstrb).
                                     .ss_tstrb (ss_tstrb).
                                     .ss_tstrb (ss_tstrb).
                                     .ss_tvalid_0 (ss_tvalid_0).
                                     .ss_tvalid_1 (ss_tvalid_1).
                                     .ss_tvalid_2 (ss_tvalid_2).
                                     .ss_tvalid_3 (ss_tvalid_3).
                                     );wire ARESET_N;
wire ASCLK;
wire [0:0] USER_PRJ_SEL;
wire a_sm_tready;
wire [pDATA_WIDTH-1:0] sm_tdata;
wire [pDATA_WIDTH-1:0] sm_tdata;
wire [pDATA_WIDTH-1:0] sm_tdata;
wire [pDATA_WIDTH-1:0] sm_tdata;
wire [2:0] sm_tid;
wire [2:0] sm_tid;
wire [2:0] sm_tid;
wire [2:0] sm_tid;
wire sm_tkeep;
wire sm_tkeep;
wire sm_tkeep;
wire sm_tkeep;
wire sm_tlast;
wire sm_tlast;
wire sm_tlast;
wire sm_tlast;
wire [3:0] sm_tstrb;
wire [3:0] sm_tstrb;
wire [3:0] sm_tstrb;
wire [3:0] sm_tstrb;
wire sm_tvalid;
wire sm_tvalid;
wire sm_tvalid;
wire sm_tvalidwire [pDATA_WIDTH-1:0] a_sm_tdata;
wire [2:0] a_sm_tid;
wire a_sm_tkeep;
wire a_sm_tlast;
wire [3:0] a_sm_tstrb;
wire a_sm_tvalid;
wire sm_tready;
wire sm_tready;
wire sm_tready;
wire sm_tready
AXIS_MSTR #(.pADDR_WIDTH(12),
            .pDATA_WIDTH(32))AXIS_MSTR (
                                     .ARESET_N (ARESET_N).
                                     .ASCLK (ASCLK).
                                     .USER_PRJ_SEL (USER_PRJ_SEL).
                                     .a_sm_tready (a_sm_tready).
                                     .sm_tdata (sm_tdata).
                                     .sm_tdata (sm_tdata).
                                     .sm_tdata (sm_tdata).
                                     .sm_tdata (sm_tdata).
                                     .sm_tid (sm_tid).
                                     .sm_tid (sm_tid).
                                     .sm_tid (sm_tid).
                                     .sm_tid (sm_tid).
                                     .sm_tkeep (sm_tkeep).
                                     .sm_tkeep (sm_tkeep).
                                     .sm_tkeep (sm_tkeep).
                                     .sm_tkeep (sm_tkeep).
                                     .sm_tlast (sm_tlast).
                                     .sm_tlast (sm_tlast).
                                     .sm_tlast (sm_tlast).
                                     .sm_tlast (sm_tlast).
                                     .sm_tstrb (sm_tstrb).
                                     .sm_tstrb (sm_tstrb).
                                     .sm_tstrb (sm_tstrb).
                                     .sm_tstrb (sm_tstrb).
                                     .sm_tvalid (sm_tvalid).
                                     .sm_tvalid (sm_tvalid).
                                     .sm_tvalid (sm_tvalid).
                                     .sm_tvalid (sm_tvalid).
                                     .a_sm_tdata (a_sm_tdata).
                                     .a_sm_tid (a_sm_tid).
                                     .a_sm_tkeep (a_sm_tkeep).
                                     .a_sm_tlast (a_sm_tlast).
                                     .a_sm_tstrb (a_sm_tstrb).
                                     .a_sm_tvalid (a_sm_tvalid).
                                     .sm_tready (sm_tready).
                                     .sm_tready (sm_tready).
                                     .sm_tready (sm_tready).
                                     .sm_tready (sm_tready).
                                     );wire ALCLK;
wire ARESET_N;
wire [0:0] USER_PRJ_SEL;
wire hi_pri_req;
wire hi_pri_req;
wire hi_pri_req;
wire hi_pri_req;
wire user_irq;
wire user_irq;
wire user_irq;
wire user_irqwire hi_pri_req;
wire user_irq
IRQ_MUX #(.pADDR_WIDTH(12),
          .pDATA_WIDTH(32))IRQ_MUX (
                                 .ALCLK (ALCLK).
                                 .ARESET_N (ARESET_N).
                                 .USER_PRJ_SEL (USER_PRJ_SEL).
                                 .hi_pri_req (hi_pri_req).
                                 .hi_pri_req (hi_pri_req).
                                 .hi_pri_req (hi_pri_req).
                                 .hi_pri_req (hi_pri_req).
                                 .user_irq (user_irq).
                                 .user_irq (user_irq).
                                 .user_irq (user_irq).
                                 .user_irq (user_irq).
                                 .hi_pri_req (hi_pri_req).
                                 .user_irq (user_irq).
                                 );wire ALCLK;
wire ARESET_N;
wire [0:0] USER_PRJ_SEL;
wire [63:0] la_data;
wire [63:0] la_data;
wire [63:0] la_data;
wire [63:0] la_datawire [63:0] la_data
LA_MUX #(.pADDR_WIDTH(12),
         .pDATA_WIDTH(32))LA_MUX (
                               .ALCLK (ALCLK).
                               .ARESET_N (ARESET_N).
                               .USER_PRJ_SEL (USER_PRJ_SEL).
                               .la_data (la_data).
                               .la_data (la_data).
                               .la_data (la_data).
                               .la_data (la_data).
                               .la_data (la_data).
                               );endmodule //USER_SUB_SYS
