module AXIL_SLAV #(parameter pADDR_WIDTH = 12,
                   parameter pDATA_WIDTH = 32)
(
	input wire ALCLK,
	input wire ARESET_N,
	input wire [0:0] USER_PRJ_SEL,
	input wire [pADDR_WIDTH-1:0] a_ls_araddr,
	input wire a_ls_arvalid,
	input wire [pADDR_WIDTH-1:0] a_ls_awaddr,
	input wire a_ls_awvalid,
	input wire [pDATA_WIDTH-1:0] a_ls_wdata,
	input wire a_ls_wstrb,
	input wire a_ls_wvalid,
	input wire a_lsrready,
	input wire arready,
	input wire arready,
	input wire arready,
	input wire arready,
	input wire awready,
	input wire awready,
	input wire awready,
	input wire awready,
	input wire [pDATA_WIDTH-1:0] rdata,
	input wire [pDATA_WIDTH-1:0] rdata,
	input wire [pDATA_WIDTH-1:0] rdata,
	input wire [pDATA_WIDTH-1:0] rdata,
	input wire rvalid,
	input wire rvalid,
	input wire rvalid,
	input wire rvalid,
	input wire wready,
	input wire wready,
	input wire wready,
	input wire wready
	output wire Arvalid_0,
	output wire [pDATA_WIDTH-1:0] Wdata,
	output wire [pDATA_WIDTH-1:0] Wdata,
	output wire [pDATA_WIDTH-1:0] Wdata,
	output wire [pDATA_WIDTH-1:0] Wdata,
	output wire a_ls_arready,
	output wire a_ls_awready,
	output wire [pDATA_WIDTH-1:0] a_ls_rdata,
	output wire a_ls_rvalid,
	output wire a_ls_wready,
	output wire [pADDR_WIDTH-1:0] araddr,
	output wire [pADDR_WIDTH-1:0] araddr,
	output wire [pADDR_WIDTH-1:0] araddr,
	output wire [pADDR_WIDTH-1:0] araddr,
	output wire arvalid_1,
	output wire arvalid_2,
	output wire arvalid_3,
	output wire [pADDR_WIDTH-1:0] awaddr,
	output wire [pADDR_WIDTH-1:0] awaddr,
	output wire [pADDR_WIDTH-1:0] awaddr,
	output wire [pADDR_WIDTH-1:0] awaddr,
	output wire awvalid_0,
	output wire awvalid_1,
	output wire awvalid_2,
	output wire awvalid_3,
	output wire rready,
	output wire rready,
	output wire rready,
	output wire rready,
	output wire wstrb_0,
	output wire wstrb_1,
	output wire wstrb_2,
	output wire wstrb_3,
	output wire wvalid_0,
	output wire wvalid_1,
	output wire wvalid_2,
	output wire wvalid_3
);

endmodule //AXIL_SLAV

